module Add32(
input [31:0] A,
input [31:0] B,
output [31:0] OUT
);
assign OUT=A+B;
endmodule
